`include "uvm_macros.svh"
import uvm_pkg::*;
`include "../../design/SPI_WRAPPER.v"
`include "SPI_Interface.sv"
`include "../Test/SPI_Seq_Item.sv"
`include "../Env/SPI_Adapter.sv"
`include "../Env/SPI_RAL.sv"
`include "../Test/SPI_Sequence.sv"
`include "../APB_Agent/APB_Sequencer.sv"
`include "../APB_Agent/APB_Driver.sv"
`include "../APB_Agent/APB_Monitor.sv"
`include "../APB_Agent/APB_Agent.sv"
`include "../SPI_Slave_agent/SPI_Slave_Sequencer.sv"
`include "../SPI_Slave_agent/SPI_Slave_Driver.sv"
`include "../SPI_Slave_agent/SPI_Slave_Monitor.sv"
`include "../SPI_Slave_agent/SPI_Slave_Agent.sv"
`include "../Env/SPI_Scoreboard.sv"
`include "../Env/Env_Config.sv"
`include "../Env/SPI_Env.sv"
`include "../Test/Test.sv"
`include "../Env/SPI_Assertions.sv"
