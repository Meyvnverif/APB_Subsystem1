class spi_coverage extends uvm_subscriber#(packet);

covergroup cg;
endgroup
endclass
